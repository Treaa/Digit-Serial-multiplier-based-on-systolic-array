`timescale 1ns / 1ps

/*
@Func: This is the testbench file for the 16 bit pipeline design of digital-serial systolic multiplier.
@Author: Jinyu Xie, Wenzhao Xie, Yuteng Huang, Hao Sun.
@Date: 2018/11/23
*/


module pipeline_16bit_tb();

parameter DATA_WIDTH = 163;
parameter B_WIDTH = 176;


reg clk;
reg rst_n;
reg [DATA_WIDTH - 1 : 0] a;
reg [DATA_WIDTH - 1 : 0] g;
reg [B_WIDTH - 1 : 0] b_total;
	
wire [DATA_WIDTH - 1 : 0] t_i_j;
reg [DATA_WIDTH - 1 : 0] t_expected;


pipeline_16bit_top tb_inst(
	.clk(clk),
	.rst_n(rst_n),
	.a(a),
	.g(g),
	.b(b_total),

	.t_i_j_out(t_i_j)
);


always begin
    clk = 1'b0;
    #10;
    clk = 1'b1;
    #10;
end

initial begin
a = 163'd0;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'd0;
t_expected = 163'd0;
rst_n = 1'b0;
#100;
rst_n = 1'b1;
#100;

a = 163'b1101100110001101100111001110110001001101000010100000000011111001110111100000110001001100011100001011001010000001110101000011000001111001000011101100011110010000010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000000111111111111111010011111010100011111110000101111111100111100110011101001110010111110000000100110101110011101111000001010101101011000100011111000110100110100111000;
t_expected = 163'b1101100000000011010001111000000011001110110001100011010000110011011010011101111100000011001000111100011111110010010010111111000000000111101010010011000101010100100;

#20;
a = 163'b0111001100101100111000110010001111111011010111101001100000111101011010100110000111110010110101101101101010101010010011001111010110010101111011111000110010001010100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000001010100101011101110000010011011011011001011011101010001110110100001000100111011001001101100000101000110100111001110101100100100110100000110001101101110000001111011;

#20;
a = 163'b0100010111010101000101110111111011011010010110011100010101100111000001110000110001111000000110110001101110100010111100100011101001010100100100111110100100110000110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000000001110010100000000101010111011010011011000001100110011000010010001010111110010110101010110100000011101101001010111100011011001011101000111110010100001011110111111;

#20;
a = 163'b0101111101100101110000001001000011100110110110010100011110100100011010100100100111000011111111101101010011001101100100001010000100101000010110111000011010110011000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000001110101001100001000110100100111111111000001101110101010011110001011111000010011000100100111000000000001000011100011001111010001010000100011101111111110001001101100;

#20;
a = 163'b1111001101001000101000110101011101000000100011010101111000001110000101110011000101011001010110011010010011110101001010000110111011000010101100111110100000101001110;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000001001111011000010100111100000101111111110110011110000011011110001101110100011011111011001101101101001010001001010111000000001000101100011110010000011000110010101101;

#20;
a = 163'b1100000111111001010101010000101001111100000010011100011001000110011110100101110011110011100011000110111111110111100110101010111000000110010110100001101100000011100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000000010100000110011011000000010101110001101101011101010001000010011101000111011010001011111101001010110011111111001010100110010001001101111011000100000011100101111111;

#20;
a = 163'b1110111101000000111000001100010001011111000001100111111010010000000000110001100101101001001010000010101010011110011001000100000111111111010100100111010010010001010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000001111110011110010011011111111011111001101110101101111000110010000111101010100111110110000010001011101011010101111100101011011101000000011111111011001100011010110000;

#20;
a = 163'b0101011110010000101111110000000111100011110000100010001111011011101001100111010001010000110011111110001010010110110001011101101000011011101111100001001100001011000;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000001000101101001001101110111111011111001111101010110011000111100110011101101101110010001111010101111100100011011000000000101100100101100111110100110001010000101110001;

#20;
a = 163'b0100000010111001010110010110111111000111110100101011101100011011110010110001000111001010111010100000000111111100011111111001011110010001010011100101100001100000100;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000000111111110101000001101011001111110101000110010110000011101000100001010111101110101000011000001110011100110001010101000011100100100101011000011001010101110010100011;

#20;
a = 163'b1110101000001100101011101011000011110001011101101011000110110001101101100111101001100000001011110100110011110101010011010101010011111101101001110011011111110010010;
g = 163'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001;
b_total = 176'b00000000000001100100101111100000000101000101111100010001100100100010110000111011011010000111011100100001111001000111000011100101101110111101001000111101101110011110101101100010;

#40;    //2 cycles(11 cycles in total)

if (t_expected == t_i_j)
	$display("1st:This data result is correct!");
else
    $display("1st:Error! The result is not as expected data.");

#20
t_expected = 163'b0101110001110001110101000111011000100111010000110111000101001000011010001111001110001011001000101100111111111011101000110001010000110101010000011011110011111010111;
if (t_expected == t_i_j)
	$display("2nd:This data result is correct!");
else
    $display("2nd:Error! The result is not as expected data.");
    
#20
t_expected = 163'b0101100110001101001010000100011001000111100101001001011011110110001100001001101111010010011010110011011001101111011000010111001000000111100100000011110000011100010;
if (t_expected == t_i_j)
	$display("3rd:This data result is correct!");
else
    $display("3rd:Error! The result is not as expected data.");
    
#20
t_expected = 163'b0000001001101111111101101110110001101010111111000000001100011111001111101011000110100001100110011001011110010100000111111110000010000100011110011000001010011101001;
if (t_expected == t_i_j)
	$display("4th:This data result is correct!");
else
    $display("4th:Error! The result is not as expected data.");
    
#20
t_expected = 163'b1110110010000111101001011111101001000100110101010111000001110010111000101101001010011110000011011110011101000111011001010011111110101011000111001010111100011001010;
if (t_expected == t_i_j)
	$display("5th:This data result is correct!");
else
    $display("5th:Error! The result is not as expected data.");
    
#20
t_expected = 163'b0100100110001100110000110110100110001110111001100001011001110100000011111101110010100100110001100100001001001001000000011011100000111111100000001010111000000101100;
if (t_expected == t_i_j)
	$display("6th:This data result is correct!");
else
    $display("6th:Error! The result is not as expected data.");
    
#20
t_expected = 163'b0111110101100010101100111110111001010000011101000010110011000010101111100011000101101010100000011001110101010011110000011100001011001001010001000110010111110110110;
if (t_expected == t_i_j)
	$display("7th:This data result is correct!");
else
    $display("7th:Error! The result is not as expected data.");

#20
t_expected = 163'b1101110101101010100010111111000011100100001101001010100000111100111110110111101001110101000001101000011110010110100101010000110101100010110001010110011000110111100;
if (t_expected == t_i_j)
	$display("8th:This data result is correct!");
else
    $display("8th:Error! The result is not as expected data.");

#20
t_expected = 163'b1010010010111101111100001001001011000100101111100001000011000011101001110101011011111111010110001010100011111101101000000100011011110001111111001011101011000010001;
if (t_expected == t_i_j)
	$display("9th:This data result is correct!");
else
    $display("9th:Error! The result is not as expected data.");

#20
t_expected = 163'b1011011001100110001110110010110010001101101001100101110110101001110110000110111100101000100010110000011110101010110001000110110001000100110001000110111101110110100;
if (t_expected == t_i_j)
	$display("10th:This data result is correct!");
else
    $display("10th:Error! The result is not as expected data.");

#10;

$finish;
end


endmodule // pipeline_16bit_tb
