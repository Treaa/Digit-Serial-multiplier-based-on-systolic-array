/*
@Func: this file is used to configure the parameter of the bit width in systolic multiplier. 
@Author: Jinyu Xie, Wenzhao Xie, Yuteng Huang, Hao Sun.
@Date: 2018/11/21
*/

`define DATA_WIDTH 163

`define N_DIGITAL 8
